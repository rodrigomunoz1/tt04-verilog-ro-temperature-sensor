`default_nettype none

(* blackbox *) module sky130_fd_sc_hd__a2111o_1(input A1, A2, B1, C1, D1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2111o_2(input A1, A2, B1, C1, D1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2111o_4(input A1, A2, B1, C1, D1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2111oi_0(input A1, A2, B1, C1, D1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2111oi_1(input A1, A2, B1, C1, D1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2111oi_2(input A1, A2, B1, C1, D1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2111oi_4(input A1, A2, B1, C1, D1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a211o_1(input A1, A2, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a211o_2(input A1, A2, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a211o_4(input A1, A2, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a211oi_1(input A1, A2, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a211oi_2(input A1, A2, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a211oi_4(input A1, A2, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21bo_1(input A1, A2, B1_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21bo_2(input A1, A2, B1_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21bo_4(input A1, A2, B1_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21boi_0(input A1, A2, B1_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21boi_1(input A1, A2, B1_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21boi_2(input A1, A2, B1_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21boi_4(input A1, A2, B1_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21o_1(input A1, A2, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21o_2(input A1, A2, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21o_4(input A1, A2, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21oi_1(input A1, A2, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21oi_2(input A1, A2, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a21oi_4(input A1, A2, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a221o_1(input A1, A2, B1, B2, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a221o_2(input A1, A2, B1, B2, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a221o_4(input A1, A2, B1, B2, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a221oi_1(input A1, A2, B1, B2, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a221oi_2(input A1, A2, B1, B2, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a221oi_4(input A1, A2, B1, B2, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a222oi_1(input A1, A2, B1, B2, C1, C2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a22o_1(input A1, A2, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a22o_2(input A1, A2, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a22o_4(input A1, A2, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a22oi_1(input A1, A2, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a22oi_2(input A1, A2, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a22oi_4(input A1, A2, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2bb2o_1(input A1_N, A2_N, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2bb2o_2(input A1_N, A2_N, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2bb2o_4(input A1_N, A2_N, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2bb2oi_1(input A1_N, A2_N, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2bb2oi_2(input A1_N, A2_N, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a2bb2oi_4(input A1_N, A2_N, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a311o_1(input A1, A2, A3, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a311o_2(input A1, A2, A3, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a311o_4(input A1, A2, A3, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a311oi_1(input A1, A2, A3, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a311oi_2(input A1, A2, A3, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a311oi_4(input A1, A2, A3, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a31o_1(input A1, A2, A3, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a31o_2(input A1, A2, A3, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a31o_4(input A1, A2, A3, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a31oi_1(input A1, A2, A3, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a31oi_2(input A1, A2, A3, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a31oi_4(input A1, A2, A3, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a32o_1(input A1, A2, A3, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a32o_2(input A1, A2, A3, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a32o_4(input A1, A2, A3, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a32oi_1(input A1, A2, A3, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a32oi_2(input A1, A2, A3, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a32oi_4(input A1, A2, A3, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a41o_1(input A1, A2, A3, A4, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a41o_2(input A1, A2, A3, A4, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a41o_4(input A1, A2, A3, A4, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__a41oi_1(input A1, A2, A3, A4, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a41oi_2(input A1, A2, A3, A4, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__a41oi_4(input A1, A2, A3, A4, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__and2_0(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and2_1(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and2_2(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and2_4(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and2b_1(input A_N, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and2b_2(input A_N, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and2b_4(input A_N, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and3_1(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and3_2(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and3_4(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and3b_1(input A_N, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and3b_2(input A_N, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and3b_4(input A_N, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4_1(input A, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4_2(input A, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4_4(input A, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4b_1(input A_N, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4b_2(input A_N, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4b_4(input A_N, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4bb_1(input A_N, B_N, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4bb_2(input A_N, B_N, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__and4bb_4(input A_N, B_N, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__buf_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__buf_12(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__buf_16(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__buf_2(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__buf_4(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__buf_6(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__buf_8(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__bufbuf_16(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__bufbuf_8(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__bufinv_16(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__bufinv_8(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkbuf_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkbuf_16(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkbuf_2(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkbuf_4(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkbuf_8(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s15_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s15_2(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s18_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s18_2(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s25_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s25_2(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s50_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkdlybuf4s50_2(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkinv_1(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkinv_16(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkinv_2(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkinv_4(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkinv_8(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkinvlp_2(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__clkinvlp_4(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__conb_1(output HI, LO); endmodule
(* blackbox *) module sky130_fd_sc_hd__decap_12(); endmodule
(* blackbox *) module sky130_fd_sc_hd__decap_3(); endmodule
(* blackbox *) module sky130_fd_sc_hd__decap_4(); endmodule
(* blackbox *) module sky130_fd_sc_hd__decap_6(); endmodule
(* blackbox *) module sky130_fd_sc_hd__decap_8(); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfbbn_1(input CLK_N, D, RESET_B, SET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfbbn_2(input CLK_N, D, RESET_B, SET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfbbp_1(input CLK, D, RESET_B, SET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfrbp_1(input CLK, D, RESET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfrbp_2(input CLK, D, RESET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfrtn_1(input CLK_N, D, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfrtp_1(input CLK, D, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfrtp_2(input CLK, D, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfrtp_4(input CLK, D, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfsbp_1(input CLK, D, SET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfsbp_2(input CLK, D, SET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfstp_1(input CLK, D, SET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfstp_2(input CLK, D, SET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfstp_4(input CLK, D, SET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfxbp_1(input CLK, D, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfxbp_2(input CLK, D, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfxtp_1(input CLK, D, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfxtp_2(input CLK, D, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dfxtp_4(input CLK, D, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__diode_2(input DIODE); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlclkp_1(input CLK, GATE, output GCLK); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlclkp_2(input CLK, GATE, output GCLK); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlclkp_4(input CLK, GATE, output GCLK); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrbn_1(input D, GATE_N, RESET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrbn_2(input D, GATE_N, RESET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrbp_1(input D, GATE, RESET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrbp_2(input D, GATE, RESET_B, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrtn_1(input D, GATE_N, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrtn_2(input D, GATE_N, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrtn_4(input D, GATE_N, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrtp_1(input D, GATE, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrtp_2(input D, GATE, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlrtp_4(input D, GATE, RESET_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlxbn_1(input D, GATE_N, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlxbn_2(input D, GATE_N, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlxbp_1(input D, GATE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlxtn_1(input D, GATE_N, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlxtn_2(input D, GATE_N, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlxtn_4(input D, GATE_N, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlxtp_1(input D, GATE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlygate4sd1_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlygate4sd2_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlygate4sd3_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlymetal6s2s_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlymetal6s4s_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__dlymetal6s6s_1(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__ebufn_1(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__ebufn_2(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__ebufn_4(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__ebufn_8(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__edfxbp_1(input CLK, D, DE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__edfxtp_1(input CLK, D, DE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvn_0(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvn_1(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvn_2(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvn_4(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvn_8(input A, TE_B, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvp_1(input A, TE, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvp_2(input A, TE, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvp_4(input A, TE, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__einvp_8(input A, TE, output Z); endmodule
(* blackbox *) module sky130_fd_sc_hd__fa_1(input A, B, CIN, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__fa_2(input A, B, CIN, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__fa_4(input A, B, CIN, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__fah_1(input A, B, CI, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__fahcin_1(input A, B, CIN, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__fahcon_1(input A, B, CI, output COUT_N, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__fill_1(); endmodule
(* blackbox *) module sky130_fd_sc_hd__fill_2(); endmodule
(* blackbox *) module sky130_fd_sc_hd__fill_4(); endmodule
(* blackbox *) module sky130_fd_sc_hd__fill_8(); endmodule
(* blackbox *) module sky130_fd_sc_hd__ha_1(input A, B, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__ha_2(input A, B, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__ha_4(input A, B, output COUT, SUM); endmodule
(* blackbox *) module sky130_fd_sc_hd__inv_1(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__inv_12(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__inv_16(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__inv_2(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__inv_4(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__inv_6(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__inv_8(input A, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_bleeder_1(input SHORT); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkbufkapwr_1(input A, KAPWR, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkbufkapwr_16(input A, KAPWR, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkbufkapwr_2(input A, KAPWR, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkbufkapwr_4(input A, KAPWR, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkbufkapwr_8(input A, KAPWR, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkinvkapwr_1(input A, KAPWR, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkinvkapwr_16(input A, KAPWR, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkinvkapwr_2(input A, KAPWR, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkinvkapwr_4(input A, KAPWR, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_clkinvkapwr_8(input A, KAPWR, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_decapkapwr_12(input KAPWR); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_decapkapwr_3(input KAPWR); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_decapkapwr_4(input KAPWR); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_decapkapwr_6(input KAPWR); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_decapkapwr_8(input KAPWR); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_inputiso0n_1(input A, SLEEP_B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_inputiso0p_1(input A, SLEEP, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_inputiso1n_1(input A, SLEEP_B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_inputiso1p_1(input A, SLEEP, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_inputisolatch_1(input D, SLEEP_B, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_isobufsrc_1(input A, SLEEP, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_isobufsrc_16(input A, SLEEP, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_isobufsrc_2(input A, SLEEP, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_isobufsrc_4(input A, SLEEP, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_isobufsrc_8(input A, SLEEP, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_isobufsrckapwr_16(input A, SLEEP, KAPWR, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1(input A, VPWRIN, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2(input A, VPWRIN, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4(input A, VPWRIN, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4(input A, output LOWLX); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1(input A, output LOWLX); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2(input A, output LOWLX); endmodule
(* blackbox *) module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4(input A, output LOWLX); endmodule
(* blackbox *) module sky130_fd_sc_hd__macro_sparecell(output LO); endmodule
(* blackbox *) module sky130_fd_sc_hd__maj3_1(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__maj3_2(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__maj3_4(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux2_1(input A0, A1, S, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux2_2(input A0, A1, S, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux2_4(input A0, A1, S, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux2_8(input A0, A1, S, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux2i_1(input A0, A1, S, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux2i_2(input A0, A1, S, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux2i_4(input A0, A1, S, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux4_1(input A0, A1, A2, A3, S0, S1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux4_2(input A0, A1, A2, A3, S0, S1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__mux4_4(input A0, A1, A2, A3, S0, S1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand2_1(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand2_2(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand2_4(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand2_8(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand2b_1(input A_N, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand2b_2(input A_N, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand2b_4(input A_N, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand3_1(input A, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand3_2(input A, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand3_4(input A, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand3b_1(input A_N, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand3b_2(input A_N, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand3b_4(input A_N, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4_1(input A, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4_2(input A, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4_4(input A, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4b_1(input A_N, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4b_2(input A_N, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4b_4(input A_N, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4bb_1(input A_N, B_N, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4bb_2(input A_N, B_N, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nand4bb_4(input A_N, B_N, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor2_1(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor2_2(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor2_4(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor2_8(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor2b_1(input A, B_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor2b_2(input A, B_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor2b_4(input A, B_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor3_1(input A, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor3_2(input A, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor3_4(input A, B, C, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor3b_1(input A, B, C_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor3b_2(input A, B, C_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor3b_4(input A, B, C_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4_1(input A, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4_2(input A, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4_4(input A, B, C, D, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4b_1(input A, B, C, D_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4b_2(input A, B, C, D_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4b_4(input A, B, C, D_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4bb_1(input A, B, C_N, D_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4bb_2(input A, B, C_N, D_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__nor4bb_4(input A, B, C_N, D_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2111a_1(input A1, A2, B1, C1, D1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2111a_2(input A1, A2, B1, C1, D1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2111a_4(input A1, A2, B1, C1, D1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2111ai_1(input A1, A2, B1, C1, D1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2111ai_2(input A1, A2, B1, C1, D1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2111ai_4(input A1, A2, B1, C1, D1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o211a_1(input A1, A2, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o211a_2(input A1, A2, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o211a_4(input A1, A2, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o211ai_1(input A1, A2, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o211ai_2(input A1, A2, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o211ai_4(input A1, A2, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21a_1(input A1, A2, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21a_2(input A1, A2, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21a_4(input A1, A2, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21ai_0(input A1, A2, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21ai_1(input A1, A2, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21ai_2(input A1, A2, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21ai_4(input A1, A2, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21ba_1(input A1, A2, B1_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21ba_2(input A1, A2, B1_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21ba_4(input A1, A2, B1_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21bai_1(input A1, A2, B1_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21bai_2(input A1, A2, B1_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o21bai_4(input A1, A2, B1_N, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o221a_1(input A1, A2, B1, B2, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o221a_2(input A1, A2, B1, B2, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o221a_4(input A1, A2, B1, B2, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o221ai_1(input A1, A2, B1, B2, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o221ai_2(input A1, A2, B1, B2, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o221ai_4(input A1, A2, B1, B2, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o22a_1(input A1, A2, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o22a_2(input A1, A2, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o22a_4(input A1, A2, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o22ai_1(input A1, A2, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o22ai_2(input A1, A2, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o22ai_4(input A1, A2, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2bb2a_1(input A1_N, A2_N, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2bb2a_2(input A1_N, A2_N, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2bb2a_4(input A1_N, A2_N, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2bb2ai_1(input A1_N, A2_N, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2bb2ai_2(input A1_N, A2_N, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o2bb2ai_4(input A1_N, A2_N, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o311a_1(input A1, A2, A3, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o311a_2(input A1, A2, A3, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o311a_4(input A1, A2, A3, B1, C1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o311ai_0(input A1, A2, A3, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o311ai_1(input A1, A2, A3, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o311ai_2(input A1, A2, A3, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o311ai_4(input A1, A2, A3, B1, C1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o31a_1(input A1, A2, A3, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o31a_2(input A1, A2, A3, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o31a_4(input A1, A2, A3, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o31ai_1(input A1, A2, A3, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o31ai_2(input A1, A2, A3, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o31ai_4(input A1, A2, A3, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o32a_1(input A1, A2, A3, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o32a_2(input A1, A2, A3, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o32a_4(input A1, A2, A3, B1, B2, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o32ai_1(input A1, A2, A3, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o32ai_2(input A1, A2, A3, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o32ai_4(input A1, A2, A3, B1, B2, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o41a_1(input A1, A2, A3, A4, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o41a_2(input A1, A2, A3, A4, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o41a_4(input A1, A2, A3, A4, B1, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__o41ai_1(input A1, A2, A3, A4, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o41ai_2(input A1, A2, A3, A4, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__o41ai_4(input A1, A2, A3, A4, B1, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__or2_0(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or2_1(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or2_2(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or2_4(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or2b_1(input A, B_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or2b_2(input A, B_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or2b_4(input A, B_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or3_1(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or3_2(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or3_4(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or3b_1(input A, B, C_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or3b_2(input A, B, C_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or3b_4(input A, B, C_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4_1(input A, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4_2(input A, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4_4(input A, B, C, D, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4b_1(input A, B, C, D_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4b_2(input A, B, C, D_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4b_4(input A, B, C, D_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4bb_1(input A, B, C_N, D_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4bb_2(input A, B, C_N, D_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__or4bb_4(input A, B, C_N, D_N, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__probe_p_8(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__probec_p_8(input A, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfbbn_1(input CLK_N, D, RESET_B, SET_B, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfbbn_2(input CLK_N, D, RESET_B, SET_B, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfbbp_1(input CLK, D, RESET_B, SET_B, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfrbp_1(input CLK, D, RESET_B, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfrbp_2(input CLK, D, RESET_B, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfrtn_1(input CLK_N, D, RESET_B, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfrtp_1(input CLK, D, RESET_B, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfrtp_2(input CLK, D, RESET_B, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfrtp_4(input CLK, D, RESET_B, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfsbp_1(input CLK, D, SET_B, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfsbp_2(input CLK, D, SET_B, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfstp_1(input CLK, D, SET_B, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfstp_2(input CLK, D, SET_B, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfstp_4(input CLK, D, SET_B, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfxbp_1(input CLK, D, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfxbp_2(input CLK, D, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfxtp_1(input CLK, D, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfxtp_2(input CLK, D, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdfxtp_4(input CLK, D, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdlclkp_1(input CLK, GATE, SCE, output GCLK); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdlclkp_2(input CLK, GATE, SCE, output GCLK); endmodule
(* blackbox *) module sky130_fd_sc_hd__sdlclkp_4(input CLK, GATE, SCE, output GCLK); endmodule
(* blackbox *) module sky130_fd_sc_hd__sedfxbp_1(input CLK, D, DE, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sedfxbp_2(input CLK, D, DE, SCD, SCE, output Q, Q_N); endmodule
(* blackbox *) module sky130_fd_sc_hd__sedfxtp_1(input CLK, D, DE, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sedfxtp_2(input CLK, D, DE, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__sedfxtp_4(input CLK, D, DE, SCD, SCE, output Q); endmodule
(* blackbox *) module sky130_fd_sc_hd__tap_1(); endmodule
(* blackbox *) module sky130_fd_sc_hd__tap_2(); endmodule
(* blackbox *) module sky130_fd_sc_hd__tapvgnd_1(); endmodule
(* blackbox *) module sky130_fd_sc_hd__tapvgnd2_1(); endmodule
(* blackbox *) module sky130_fd_sc_hd__tapvpwrvgnd_1(); endmodule
(* blackbox *) module sky130_fd_sc_hd__xnor2_1(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__xnor2_2(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__xnor2_4(input A, B, output Y); endmodule
(* blackbox *) module sky130_fd_sc_hd__xnor3_1(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xnor3_2(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xnor3_4(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xor2_1(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xor2_2(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xor2_4(input A, B, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xor3_1(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xor3_2(input A, B, C, output X); endmodule
(* blackbox *) module sky130_fd_sc_hd__xor3_4(input A, B, C, output X); endmodule
